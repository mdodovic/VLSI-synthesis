module hex (
	input [3:0] in,
	output reg [6:0] out
);

/*
 *                              A
 *                           *******
 *                         *         *
 *                       F *         * B
 *                         *    G    *
 *                           *******
 *                         *         *
 *                       E *         * C
 *                         *    D    *
 *                           *******
 * 
 * 1 means light
 * It should be inverted (~) on assgin!
 * |-----|||-----|-----|-----|-----|-----|-----|-----|||-----|
 * | DIG |||  G  |  F  |  E  |  D  |  C  |  B  |  A  ||| VAL |
 * |-----|||-----|-----|-----|-----|-----|-----|-----|||-----|
 * |  0  |||  0  |  1  |  1  |  1  |  1  |  1  |  1  ||| 3F  | 
 * |  1  |||  0  |  0  |  0  |  0  |  1  |  1  |  0  ||| 06  | 
 * |  2  |||  1  |  0  |  1  |  1  |  0  |  0  |  0  ||| 58  | 
 * |  3  |||  1  |  0  |  0  |  1  |  1  |  1  |  1  ||| 4F  |
 * |  4  |||  1  |  1  |  0  |  0  |  1  |  1  |  0  ||| 66  |
 * |  5  |||  1  |  1  |  0  |  1  |  1  |  0  |  1  ||| 6D  |
 * |  6  |||  1  |  1  |  1  |  1  |  1  |  0  |  1  ||| 7D  |
 * |  7  |||  0  |  0  |  0  |  0  |  1  |  1  |  1  ||| 07  |
 * |  8  |||  1  |  1  |  1  |  1  |  1  |  1  |  1  ||| 7F  |
 * |  9  |||  1  |  0  |  1  |  1  |  1  |  1  |  1  ||| 6F  |
 * |  A  |||  1  |  1  |  1  |  0  |  1  |  1  |  1  ||| 77  |
 * |  b  |||  1  |  1  |  1  |  1  |  1  |  0  |  0  ||| 7C  | 
 * |  C  |||  0  |  1  |  1  |  1  |  0  |  0  |  1  ||| 39  | 
 * |  d  |||  1  |  0  |  1  |  1  |  1  |  1  |  0  ||| 5E  | 
 * |  E  |||  1  |  1  |  1  |  1  |  0  |  0  |  1  ||| 79  |
 * |  F  |||  1  |  1  |  1  |  0  |  0  |  0  |  1  ||| 71  |
 * |-----|||-----|-----|-----|-----|-----|-----|-----|||-----|
 *
 */

	always @(*) begin
        case (in)
            4'b0000: out = ~7'h3F; // 7seg is active in logic zero 
            4'b0001: out = ~7'h06;  
            4'b0010: out = ~7'h5B;  
            4'b0011: out = ~7'h4F;
            4'b0100: out = ~7'h66;
            4'b0101: out = ~7'h6D;
            4'b0110: out = ~7'h7D;
            4'b0111: out = ~7'h07;
            4'b1000: out = ~7'h7F;
            4'b1001: out = ~7'h6F;
            4'b1010: out = ~7'h77;
            4'b1011: out = ~7'h7C;
            4'b1100: out = ~7'h39;
            4'b1101: out = ~7'h5E;
            4'b1110: out = ~7'h79;
            4'b1111: out = ~7'h71;
        endcase
	end
	
endmodule